module top(
	input  clk,
	input  [7:0]address,
	input  sw,
	input  [3:0]ch,
	output [3:0]anode,
	output [7:0]segment
);

endmodule